VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ExampleDCO
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN ExampleDCO 0 0 ;
  SIZE 123.936 BY 125.536 ;
  SYMMETRY X Y ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT 
      LAYER M5 ;
        RECT 3.024 121.536 3.8 125.536 ;
    END 
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT 
      LAYER M5 ;
        RECT 1.728 121.536 2.5 125.536 ;
    END 
  END VSS
  PIN dither
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.384 1.2 0.768 ;
    END 
  END dither
  PIN row_sel_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.536 1.2 1.92 ;
    END 
  END row_sel_b[0]
  PIN row_sel_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.688 1.2 3.072 ;
    END 
  END row_sel_b[1]
  PIN row_sel_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.84 1.2 4.224 ;
    END 
  END row_sel_b[2]
  PIN row_sel_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.992 1.2 5.376 ;
    END 
  END row_sel_b[3]
  PIN row_sel_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.144 1.2 6.528 ;
    END 
  END row_sel_b[4]
  PIN row_sel_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.296 1.2 7.68 ;
    END 
  END row_sel_b[5]
  PIN row_sel_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.448 1.2 8.832 ;
    END 
  END row_sel_b[6]
  PIN row_sel_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.6 1.2 9.984 ;
    END 
  END row_sel_b[7]
  PIN row_sel_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.752 1.2 11.136 ;
    END 
  END row_sel_b[8]
  PIN row_sel_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.904 1.2 12.288 ;
    END 
  END row_sel_b[9]
  PIN row_sel_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.056 1.2 13.44 ;
    END 
  END row_sel_b[10]
  PIN row_sel_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.208 1.2 14.592 ;
    END 
  END row_sel_b[11]
  PIN row_sel_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.36 1.2 15.744 ;
    END 
  END row_sel_b[12]
  PIN row_sel_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.512 1.2 16.896 ;
    END 
  END row_sel_b[13]
  PIN row_sel_b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.664 1.2 18.048 ;
    END 
  END row_sel_b[14]
  PIN row_sel_b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.816 1.2 19.2 ;
    END 
  END row_sel_b[15]
  PIN col_sel_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.968 1.2 20.352 ;
    END 
  END col_sel_b[0]
  PIN col_sel_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.12 1.2 21.504 ;
    END 
  END col_sel_b[1]
  PIN col_sel_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 22.272 1.2 22.656 ;
    END 
  END col_sel_b[2]
  PIN col_sel_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.424 1.2 23.808 ;
    END 
  END col_sel_b[3]
  PIN col_sel_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.576 1.2 24.96 ;
    END 
  END col_sel_b[4]
  PIN col_sel_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.728 1.2 26.112 ;
    END 
  END col_sel_b[5]
  PIN col_sel_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 26.88 1.2 27.264 ;
    END 
  END col_sel_b[6]
  PIN col_sel_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 28.032 1.2 28.416 ;
    END 
  END col_sel_b[7]
  PIN col_sel_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 29.184 1.2 29.568 ;
    END 
  END col_sel_b[8]
  PIN col_sel_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 30.336 1.2 30.72 ;
    END 
  END col_sel_b[9]
  PIN col_sel_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.488 1.2 31.872 ;
    END 
  END col_sel_b[10]
  PIN col_sel_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 32.64 1.2 33.024 ;
    END 
  END col_sel_b[11]
  PIN col_sel_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 33.792 1.2 34.176 ;
    END 
  END col_sel_b[12]
  PIN col_sel_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 34.944 1.2 35.328 ;
    END 
  END col_sel_b[13]
  PIN code_regulator[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 36.096 1.2 36.48 ;
    END 
  END code_regulator[0]
  PIN code_regulator[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 37.248 1.2 37.632 ;
    END 
  END code_regulator[1]
  PIN code_regulator[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 38.4 1.2 38.784 ;
    END 
  END code_regulator[2]
  PIN code_regulator[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 39.552 1.2 39.936 ;
    END 
  END code_regulator[3]
  PIN code_regulator[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 40.704 1.2 41.088 ;
    END 
  END code_regulator[4]
  PIN code_regulator[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 41.856 1.2 42.24 ;
    END 
  END code_regulator[5]
  PIN code_regulator[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 43.008 1.2 43.392 ;
    END 
  END code_regulator[6]
  PIN code_regulator[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 44.16 1.2 44.544 ;
    END 
  END code_regulator[7]
  PIN sleep_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 45.312 1.2 45.696 ;
    END 
  END sleep_b
  PIN clock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 122.736 0.384 123.936 0.768 ;
    END 
  END clock
  OBS 
    LAYER M1 ;
      RECT 1.2 0.0 122.736 121.536 ;
    LAYER M2 ;
      RECT 1.2 0.0 122.736 121.536 ;
    LAYER M3 ;
      RECT 1.2 0.0 122.736 121.536 ;
    LAYER M4 ;
      RECT 1.2 0.0 122.736 121.536 ;
    LAYER M5 ;
      RECT 1.2 0.0 122.736 121.536 ;
    LAYER M6 ;
      RECT 1.2 0.0 122.736 121.536 ;
    LAYER M7 ;
      RECT 1.2 0.0 122.736 121.536 ;
    LAYER M8 ;
      RECT 1.2 0.0 122.736 121.536 ;
    LAYER M9 ;
      RECT 1.2 0.0 122.736 121.536 ;
  END 
END ExampleDCO

END LIBRARY
