VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ExampleDCO
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN ExampleDCO 0 0 ;
  SIZE 129.536 BY 125.536 ;
  SYMMETRY X Y ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT 
      LAYER M5 ;
        RECT 10.608 121.536 11.088 125.536 ;
    END 
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT 
      LAYER M5 ;
        RECT 11.712 121.536 12.192 125.536 ;
    END 
  END VSS
  PIN dither
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.384 4.0 0.768 ;
    END 
  END dither
  PIN row_sel_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.536 4.0 1.92 ;
    END 
  END row_sel_b[0]
  PIN row_sel_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.688 4.0 3.072 ;
    END 
  END row_sel_b[1]
  PIN row_sel_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.84 4.0 4.224 ;
    END 
  END row_sel_b[2]
  PIN row_sel_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.992 4.0 5.376 ;
    END 
  END row_sel_b[3]
  PIN row_sel_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.144 4.0 6.528 ;
    END 
  END row_sel_b[4]
  PIN row_sel_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.296 4.0 7.68 ;
    END 
  END row_sel_b[5]
  PIN row_sel_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.448 4.0 8.832 ;
    END 
  END row_sel_b[6]
  PIN row_sel_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.6 4.0 9.984 ;
    END 
  END row_sel_b[7]
  PIN row_sel_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.752 4.0 11.136 ;
    END 
  END row_sel_b[8]
  PIN row_sel_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.904 4.0 12.288 ;
    END 
  END row_sel_b[9]
  PIN row_sel_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.056 4.0 13.44 ;
    END 
  END row_sel_b[10]
  PIN row_sel_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.208 4.0 14.592 ;
    END 
  END row_sel_b[11]
  PIN row_sel_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.36 4.0 15.744 ;
    END 
  END row_sel_b[12]
  PIN row_sel_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.512 4.0 16.896 ;
    END 
  END row_sel_b[13]
  PIN row_sel_b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.664 4.0 18.048 ;
    END 
  END row_sel_b[14]
  PIN row_sel_b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.816 4.0 19.2 ;
    END 
  END row_sel_b[15]
  PIN col_sel_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.968 4.0 20.352 ;
    END 
  END col_sel_b[0]
  PIN col_sel_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.12 4.0 21.504 ;
    END 
  END col_sel_b[1]
  PIN col_sel_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 22.272 4.0 22.656 ;
    END 
  END col_sel_b[2]
  PIN col_sel_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.424 4.0 23.808 ;
    END 
  END col_sel_b[3]
  PIN col_sel_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.576 4.0 24.96 ;
    END 
  END col_sel_b[4]
  PIN col_sel_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.728 4.0 26.112 ;
    END 
  END col_sel_b[5]
  PIN col_sel_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 26.88 4.0 27.264 ;
    END 
  END col_sel_b[6]
  PIN col_sel_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 28.032 4.0 28.416 ;
    END 
  END col_sel_b[7]
  PIN col_sel_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 29.184 4.0 29.568 ;
    END 
  END col_sel_b[8]
  PIN col_sel_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 30.336 4.0 30.72 ;
    END 
  END col_sel_b[9]
  PIN col_sel_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.488 4.0 31.872 ;
    END 
  END col_sel_b[10]
  PIN col_sel_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 32.64 4.0 33.024 ;
    END 
  END col_sel_b[11]
  PIN col_sel_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 33.792 4.0 34.176 ;
    END 
  END col_sel_b[12]
  PIN col_sel_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 34.944 4.0 35.328 ;
    END 
  END col_sel_b[13]
  PIN code_regulator[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 36.096 4.0 36.48 ;
    END 
  END code_regulator[0]
  PIN code_regulator[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 37.248 4.0 37.632 ;
    END 
  END code_regulator[1]
  PIN code_regulator[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 38.4 4.0 38.784 ;
    END 
  END code_regulator[2]
  PIN code_regulator[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 39.552 4.0 39.936 ;
    END 
  END code_regulator[3]
  PIN code_regulator[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 40.704 4.0 41.088 ;
    END 
  END code_regulator[4]
  PIN code_regulator[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 41.856 4.0 42.24 ;
    END 
  END code_regulator[5]
  PIN code_regulator[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 43.008 4.0 43.392 ;
    END 
  END code_regulator[6]
  PIN code_regulator[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 44.16 4.0 44.544 ;
    END 
  END code_regulator[7]
  PIN sleep_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 45.312 4.0 45.696 ;
    END 
  END sleep_b
  PIN clock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 125.536 0.384 129.536 0.768 ;
    END 
  END clock
  OBS 
    LAYER M1 ;
      RECT 4.0 0.0 125.536 121.536 ;
    LAYER M2 ;
      RECT 4.0 0.0 125.536 121.536 ;
    LAYER M3 ;
      RECT 4.0 0.0 125.536 121.536 ;
    LAYER M4 ;
      RECT 4.0 0.0 125.536 121.536 ;
    LAYER M5 ;
      RECT 4.0 0.0 125.536 121.536 ;
    LAYER M6 ;
      RECT 4.0 0.0 125.536 121.536 ;
    LAYER M7 ;
      RECT 4.0 0.0 125.536 121.536 ;
    LAYER M8 ;
      RECT 0.0 0.0 129.536 121.536 ;
    LAYER M9 ;
      RECT 0.0 0.0 129.536 121.536 ;
    LAYER Pad ;
      RECT 0.0 0.0 129.536 121.536 ;
  END 
END ExampleDCO

END LIBRARY
