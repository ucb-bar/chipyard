module ExampleVerilogTLDevice #(
                                parameter CTRL_ADDR_BITS,
                                parameter CTRL_DATA_BITS,
                                parameter CTRL_SOURCE_BITS,
                                parameter CTRL_SINK_BITS,
                                parameter CTRL_SIZE_BITS,
                                parameter CLIENT_ADDR_BITS,
                                parameter CLIENT_DATA_BITS,
                                parameter CLIENT_SOURCE_BITS,
                                parameter CLIENT_SINK_BITS,
                                parameter CLIENT_SIZE_BITS
                                )(
  input                             tl_client_a_ready,
  output                            tl_client_a_valid,
  output [2:0]                      tl_client_a_bits_opcode,
  output [2:0]                      tl_client_a_bits_param,
  output [CLIENT_SIZE_BITS-1:0]     tl_client_a_bits_size,
  output [CLIENT_SOURCE_BITS-1:0]   tl_client_a_bits_source,
  output [CLIENT_ADDR_BITS-1:0]     tl_client_a_bits_address,
  output [(CLIENT_DATA_BITS/8)-1:0] tl_client_a_bits_mask,
  output [CLIENT_DATA_BITS-1:0]     tl_client_a_bits_data,
  output                            tl_client_a_bits_corrupt,
  output                            tl_client_d_ready,
  input                             tl_client_d_valid,
  input [2:0]                       tl_client_d_bits_opcode,
  input [1:0]                       tl_client_d_bits_param,
  input [CLIENT_SIZE_BITS-1:0]      tl_client_d_bits_size,
  input [CLIENT_SOURCE_BITS-1:0]    tl_client_d_bits_source,
  input [CLIENT_SINK_BITS-1:0]      tl_client_d_bits_sink,
  input                             tl_client_d_bits_denied,
  input [CLIENT_DATA_BITS-1:0]      tl_client_d_bits_data,
  input                             tl_client_d_bits_corrupt,
  output                            tl_ctrl_a_ready,
  input                             tl_ctrl_a_valid,
  input [2:0]                       tl_ctrl_a_bits_opcode,
  input [2:0]                       tl_ctrl_a_bits_param,
  input [CTRL_SIZE_BITS-1:0]        tl_ctrl_a_bits_size,
  input [CTRL_SOURCE_BITS-1:0]      tl_ctrl_a_bits_source,
  input [CTRL_ADDR_BITS-1:0]        tl_ctrl_a_bits_address,
  input [(CTRL_DATA_BITS/8)-1:0]    tl_ctrl_a_bits_mask,
  input [CTRL_DATA_BITS-1:0]        tl_ctrl_a_bits_data,
  input                             tl_ctrl_a_bits_corrupt,
  input                             tl_ctrl_d_ready,
  output                            tl_ctrl_d_valid,
  output [2:0]                      tl_ctrl_d_bits_opcode,
  output [1:0]                      tl_ctrl_d_bits_param,
  output [CTRL_SIZE_BITS-1:0]       tl_ctrl_d_bits_size,
  output [CTRL_SOURCE_BITS-1:0]     tl_ctrl_d_bits_source,
  output [CTRL_SINK_BITS-1:0]       tl_ctrl_d_bits_sink,
  output                            tl_ctrl_d_bits_denied,
  output [CTRL_DATA_BITS-1:0]       tl_ctrl_d_bits_data,
  output                            tl_ctrl_d_bits_corrupt,
  input                             clock,
  input                             reset
);

endmodule
