VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ExampleDCO
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN ExampleDCO 0 0 ;
  SIZE 128.0 BY 128.0 ;
  SYMMETRY X Y ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M7 ;
        RECT 32.96 124.0 33.6 128.0 ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 93.12 124.0 93.76 128.0 ; 
    END
  END VSS
  PIN col_sel_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 113.28 4.0 113.664 ; 
    END
  END col_sel_b[13]
  PIN col_sel_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 107.648 4.0 108.032 ; 
    END
  END col_sel_b[11]
  PIN col_sel_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 90.752 4.0 91.136 ; 
    END
  END col_sel_b[5]
  PIN col_sel_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 110.464 4.0 110.848 ; 
    END
  END col_sel_b[12]
  PIN col_sel_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 104.832 4.0 105.216 ; 
    END
  END col_sel_b[10]
  PIN col_sel_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 102.016 4.0 102.4 ; 
    END
  END col_sel_b[9]
  PIN col_sel_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 99.2 4.0 99.584 ; 
    END
  END col_sel_b[8]
  PIN col_sel_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 96.384 4.0 96.768 ; 
    END
  END col_sel_b[7]
  PIN col_sel_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 93.568 4.0 93.952 ; 
    END
  END col_sel_b[6]
  PIN col_sel_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 87.936 4.0 88.32 ; 
    END
  END col_sel_b[4]
  PIN col_sel_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 85.12 4.0 85.504 ; 
    END
  END col_sel_b[3]
  PIN col_sel_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 82.304 4.0 82.688 ; 
    END
  END col_sel_b[2]
  PIN col_sel_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 79.488 4.0 79.872 ; 
    END
  END col_sel_b[1]
  PIN col_sel_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 76.672 4.0 77.056 ; 
    END
  END col_sel_b[0]
  PIN row_sel_b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 71.04 4.0 71.424 ; 
    END
  END row_sel_b[14]
  PIN row_sel_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 68.224 4.0 68.608 ; 
    END
  END row_sel_b[13]
  PIN row_sel_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 65.408 4.0 65.792 ; 
    END
  END row_sel_b[12]
  PIN row_sel_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 62.592 4.0 62.976 ; 
    END
  END row_sel_b[11]
  PIN row_sel_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 59.776 4.0 60.16 ; 
    END
  END row_sel_b[10]
  PIN row_sel_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 56.96 4.0 57.344 ; 
    END
  END row_sel_b[9]
  PIN row_sel_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 54.144 4.0 54.528 ; 
    END
  END row_sel_b[8]
  PIN row_sel_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 51.328 4.0 51.712 ; 
    END
  END row_sel_b[7]
  PIN row_sel_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 48.512 4.0 48.896 ; 
    END
  END row_sel_b[6]
  PIN row_sel_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 45.696 4.0 46.08 ; 
    END
  END row_sel_b[5]
  PIN row_sel_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 42.88 4.0 43.264 ; 
    END
  END row_sel_b[4]
  PIN row_sel_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 40.064 4.0 40.448 ; 
    END
  END row_sel_b[3]
  PIN row_sel_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 37.248 4.0 37.632 ; 
    END
  END row_sel_b[2]
  PIN row_sel_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 34.432 4.0 34.816 ; 
    END
  END row_sel_b[1]
  PIN row_sel_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 31.616 4.0 32.0 ; 
    END
  END row_sel_b[0]
  PIN code_regulator[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 28.8 4.0 29.184 ; 
    END
  END code_regulator[7]
  PIN code_regulator[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 25.984 4.0 26.368 ; 
    END
  END code_regulator[6]
  PIN code_regulator[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 23.168 4.0 23.552 ; 
    END
  END code_regulator[5]
  PIN code_regulator[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 20.352 4.0 20.736 ; 
    END
  END code_regulator[4]
  PIN code_regulator[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 17.536 4.0 17.92 ; 
    END
  END code_regulator[3]
  PIN code_regulator[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 14.72 4.0 15.104 ; 
    END
  END code_regulator[2]
  PIN code_regulator[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 11.904 4.0 12.288 ; 
    END
  END code_regulator[1]
  PIN code_regulator[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 9.088 4.0 9.472 ; 
    END
  END code_regulator[0]
  PIN row_sel_b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 73.856 4.0 74.24 ; 
    END
  END row_sel_b[15]
  PIN dither
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 6.272 4.0 6.656 ; 
    END
  END dither
  PIN sleep_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.792 0.0 10.176 4.0 ; 
    END
  END sleep_b
  PIN clock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 124.0 70.864 128.0 71.248 ; 
    END
  END clock
  OBS
    LAYER M1 ;
      RECT 4.0 4.0 124.0 124.0 ; 
    LAYER M2 ;
      RECT 4.0 4.0 124.0 124.0 ; 
    LAYER M3 ;
      RECT 4.0 4.0 124.0 124.0 ; 
    LAYER M4 ;
      RECT 4.0 4.0 124.0 124.0 ; 
    LAYER M5 ;
      RECT 4.0 4.0 124.0 124.0 ;
    LAYER M6 ;
      RECT 4.0 4.0 124.0 124.0 ; 
    LAYER M7 ;
      RECT 4.0 4.0 124.0 124.0 ; 
    LAYER M8 ;
      RECT 0.0 0.0 128.0 128.0 ; 
    LAYER M9 ;
      RECT 0.0 0.0 128.0 128.0 ; 
    LAYER Pad ;
      RECT 0.0 0.0 128.0 128.0 ; 
  END
END ExampleDCO

END LIBRARY
