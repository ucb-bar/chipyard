VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ExampleDCO
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ExampleDCO 0 0 ;
  SIZE 32.001 BY 32 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
        RECT 8.24 31 8.4 32 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
        RECT 23.28 31 23.44 32 ;
    END
  END VSS
  PIN col_sel_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 28.32 1 28.416 ;
    END
  END col_sel_b[13]
  PIN col_sel_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 26.912 1 27.008 ;
    END
  END col_sel_b[11]
  PIN col_sel_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 22.688 1 22.784 ;
    END
  END col_sel_b[5]
  PIN col_sel_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 27.616 1 27.712 ;
    END
  END col_sel_b[12]
  PIN col_sel_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 26.208 1 26.304 ;
    END
  END col_sel_b[10]
  PIN col_sel_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 25.504 1 25.6 ;
    END
  END col_sel_b[9]
  PIN col_sel_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 24.8 1 24.896 ;
    END
  END col_sel_b[8]
  PIN col_sel_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 24.096 1 24.192 ;
    END
  END col_sel_b[7]
  PIN col_sel_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 23.392 1 23.488 ;
    END
  END col_sel_b[6]
  PIN col_sel_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 21.984 1 22.08 ;
    END
  END col_sel_b[4]
  PIN col_sel_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 21.28 1 21.376 ;
    END
  END col_sel_b[3]
  PIN col_sel_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 20.576 1 20.672 ;
    END
  END col_sel_b[2]
  PIN col_sel_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 19.872 1 19.968 ;
    END
  END col_sel_b[1]
  PIN col_sel_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 19.168 1 19.264 ;
    END
  END col_sel_b[0]
  PIN row_sel_b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 17.76 1 17.856 ;
    END
  END row_sel_b[14]
  PIN row_sel_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 17.056 1 17.152 ;
    END
  END row_sel_b[13]
  PIN row_sel_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 16.352 1 16.448 ;
    END
  END row_sel_b[12]
  PIN row_sel_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 15.648 1 15.744 ;
    END
  END row_sel_b[11]
  PIN row_sel_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 14.944 1 15.04 ;
    END
  END row_sel_b[10]
  PIN row_sel_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 14.24 1 14.336 ;
    END
  END row_sel_b[9]
  PIN row_sel_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 13.536 1 13.632 ;
    END
  END row_sel_b[8]
  PIN row_sel_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 12.832 1 12.928 ;
    END
  END row_sel_b[7]
  PIN row_sel_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 12.128 1 12.224 ;
    END
  END row_sel_b[6]
  PIN row_sel_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 11.424 1 11.52 ;
    END
  END row_sel_b[5]
  PIN row_sel_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 10.72 1 10.816 ;
    END
  END row_sel_b[4]
  PIN row_sel_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 10.016 1 10.112 ;
    END
  END row_sel_b[3]
  PIN row_sel_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 9.312 1 9.408 ;
    END
  END row_sel_b[2]
  PIN row_sel_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 8.608 1 8.704 ;
    END
  END row_sel_b[1]
  PIN row_sel_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 7.904 1 8 ;
    END
  END row_sel_b[0]
  PIN code_regulator[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 7.2 1 7.296 ;
    END
  END code_regulator[7]
  PIN code_regulator[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 6.496 1 6.592 ;
    END
  END code_regulator[6]
  PIN code_regulator[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 5.792 1 5.888 ;
    END
  END code_regulator[5]
  PIN code_regulator[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 5.088 1 5.184 ;
    END
  END code_regulator[4]
  PIN code_regulator[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 4.384 1 4.48 ;
    END
  END code_regulator[3]
  PIN code_regulator[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 3.68 1 3.776 ;
    END
  END code_regulator[2]
  PIN code_regulator[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 2.976 1 3.072 ;
    END
  END code_regulator[1]
  PIN code_regulator[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 2.272 1 2.368 ;
    END
  END code_regulator[0]
  PIN row_sel_b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 18.464 1 18.56 ;
    END
  END row_sel_b[15]
  PIN dither
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 1.568 1 1.664 ;
    END
  END dither
  PIN sleep_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.448 0 2.544 1 ;
    END
  END sleep_b
  PIN clock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31 17.716 32 17.812 ;
    END
  END clock
  OBS
    LAYER M1 ;
      RECT 1 1 31 31 ;
    LAYER M2 ;
      RECT 1 1 31 31 ;
    LAYER M3 ;
      RECT 1 1 31 31 ;
    LAYER M4 ;
      RECT 1 1 31 31 ;
    LAYER M6 ;
      RECT 1 1 31 31 ;
    LAYER M7 ;
      RECT 1 1 31 31 ;
    LAYER M8 ;
      RECT 1 1 31 31 ;
    LAYER M9 ;
      RECT 1 1 31 31 ;
  END
END ExampleDCO

END LIBRARY
